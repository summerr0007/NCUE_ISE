module rain();

endmodule;